module cnn (
    input w_data[31:0];
    input addr[1:0];
    output r_data[31:0];
)

 sram dut(

 );


endmodule


module sram()

endmodule